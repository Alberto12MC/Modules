-------------------------------------------------------
--! @file  fsm.vhd
--! @brief
--! @todo
--! @defgroup fsm
-------------------------------------------------------

--! Standard library.
library ieee;
--! Logic elements.
use ieee.std_logic_1164.all;
--! arithmetic functions.
use ieee.numeric_std.all;

--! @brief   implementation
--! @details implementation of xxx
--! @ingroup fsm

entity fsm is
  generic(

  );
  port (
         -- Common
         clk   : in std_logic;
         reset : in std_logic;
  );
end fsm;

architecture rtl of fsm is


begin


end rtl;
